`timescale 1ns / 1ps

///////////////////////////////////////////////////////////////////

//GROUP NUMBER  - A05
//GROUP MEMBERS - ASHNA JAIN(201501008)
//					 - CHARMI CHOKSHI(201501021)
//              - MANASI DUBEY(201501051)
//DESCRIPTION:  - This is the Register Bank block of microprocessor.

///////////////////////////////////////////////////////////////////


module register_bank_module(ins, RW_dm, ans_ex, mux_ans_dm, ans_wb, imm, mux_sel_A, mux_sel_B, imm_sel, clk, reset, A, B);

output [7:0] A, B;		//initializing outputs which are of 8 bits

input [19:0] ins;			//initializing input which are of 20 bits
input [4:0] RW_dm;		//initializing input which are of 5 bits
input [7:0] ans_ex, mux_ans_dm, ans_wb, imm;			//initializing input which are of 8 bits
input [1:0] mux_sel_A, mux_sel_B;		//initializing input which are of 2 bits
input imm_sel, clk, reset;			//initializing input which are of 1 bits

wire [4:0] RA, RB;			//initializing wire which are of 5 bits
reg [7:0] reg_A, reg_B;			//initializing registers which are of 8 bits
wire [7:0] temp_B;			//initializing wires which are of 8 bits
reg [7:0] arr[0:31];		//initializing register which are of 8 bits and allocating such 32 addresses to it
wire [7:0] arr_t,reg_A_t,reg_B_t;

assign RA = ins[9:5];		//assigning bits from 9 to 5 of ins to RA
assign RB = ins[4:0];		//assignning the first 5 bits of ins to RB

initial 
begin

	arr[0] <= 0;			//using non blocking approch giving the value 0(data) to a[0](Location) to Initialize Reg Bank
	arr[1] <= 1;			//countinuing for 32 bits
	arr[2] <= 2;
	arr[3] <= 3;
	arr[4] <= 4;
	arr[5] <= 5;
	arr[6] <= 6;
	arr[7] <= 7;
	arr[8] <= 8;
	arr[9] <= 9;
	arr[10] <= 10;
	arr[11] <= 11;
	arr[12] <= 12;
	arr[13] <= 13;
	arr[14] <= 14;
	arr[15] <= 15;
	arr[16] <= 16;
	arr[17] <= 17;
	arr[18] <= 18;
	arr[19] <= 19;
	arr[20] <= 20;
	arr[21] <= 21;
	arr[22] <= 22;
	arr[23] <= 23;
	arr[24] <= 24;
	arr[25] <= 25;
	arr[26] <= 26;
	arr[27] <= 27;
	arr[28] <= 28;
	arr[29] <= 29;
	arr[30] <= 30;
	arr[31] <= 31;
	
end

assign arr_t = (reset==1'b1) ? mux_ans_dm : 8'b00000000;		//assigning mux_ans_dm to arr_t when reset is 1 else 0 (arr_t is a wire that gives the value to arr[RW_dm] at posedge clk)
assign reg_A_t= (reset==1'b1) ? arr[RA] : 8'b00000000;		//assigning arr[RA] to reg_A_t when reset is 1 else 0 (reg_A_t is a wire that gives the value to reg_A at posedge clk)
assign reg_B_t= (reset==1'b1) ? arr[RB] : 8'b00000000;		//assigning arr[RB] to reg_B_t when reset is 1 else 0 (reg_B_t is a wire that gives the value to reg_B at posedge clk)

always@(posedge clk)			//this block will execute whene the clock is at posedge
begin
  		arr[RW_dm] <= arr_t;		//assigning the value of  arr_t to arr[RW_dm] at the address RW_dm
      reg_A <= reg_A_t;			//assignning the value of reg_A_t to reg_A
		reg_B <= reg_B_t;			//assignning the value of reg_B_t to reg_B
end


/*		according to signals generated by dependency check block(mux_sel_A and mux_sel_B),
		assigning the value to outputs A and B from ans_wb, ans_ex, mux_ans_dm, reg_A/reg_B
		
		if any immidiate number is given than taking that number as output B
*/

assign A = (mux_sel_A == 2'b00 ?reg_A:(mux_sel_A == 2'b01 ?ans_ex:(mux_sel_A == 2'b10 ?mux_ans_dm:(mux_sel_A == 2'b11 ?ans_wb:8'b00000000))));		//creating MUX using ternanry operator
assign temp_B = (mux_sel_B == 2'b00 ?reg_B:(mux_sel_B == 2'b01 ?ans_ex:(mux_sel_B == 2'b10 ?mux_ans_dm:(mux_sel_B == 2'b11 ?ans_wb:8'b00000000))));		//creating MUX using ternanry operator
assign B = (imm_sel == 1'b0 ?temp_B:(imm_sel == 1'b1 ?imm:8'b00000000));			//creating MUX using ternanry operator

endmodule		//body of code ends here