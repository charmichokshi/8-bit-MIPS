`timescale 1ns / 1ps

///////////////////////////////////////////////////////////////////

//GROUP NUMBER  - A05
//GROUP MEMBERS - ASHNA JAIN(201501008)
//					 - CHARMI CHOKSHI(201501021)
//              - MANASI DUBEY(201501051)
//DESCRIPTION:  - This is the Execution block of microprocessor.

///////////////////////////////////////////////////////////////////
module execution_module(flag_ex,ans_ex,data_out,B_Bypass,mem_en_ex,mem_rw_ex,mem_mux_sel_ex,RW_ex,A,B,data_in,op_dec,clk,mem_en_dec,mem_rw_dec,mem_mux_sel_dec,RW_dec,reset);

//output declaration
output [3:0] flag_ex;
output reg [7:0] ans_ex;
output reg [7:0] data_out,B_Bypass;
output reg mem_en_ex,mem_rw_ex,mem_mux_sel_ex;
output reg [4:0] RW_ex;

//input declaration
input [7:0] A,B,data_in;
input [4:0] op_dec;
input [4:0] RW_dec;
input clk,reset;
input mem_en_dec,mem_rw_dec,mem_mux_sel_dec;

//wire declaration
wire [7:0] a1,a2,a4,a5,a6,a7,a22,a23,a24,c1,ans_temp;
wire flag_temp,t1,t2,t3,t4,t5,t6,carry1,carry2,flag1,flag2,flag3,flag4,carry;

wire r1,r2,r3,r4;
wire [7:0] data_out_buff;
wire [7:0] ans_ex_t, data_out_t, B_Bypass_t;
wire mem_en_ex_t, mem_rw_ex_t, mem_mux_sel_ex_t;
wire [4:0] RW_ex_t;

//This block calculates the sum of A and B and stores the carry in carry1 
assign {carry1,a1}=A[7:0]+ B[7:0];	//finding the sum of A and B, storing the sum in a1 and carry in carry1
assign {flag1}=A[5:0]+B[5:0];		//calculating the sum of first six bits and storing the carry generated by adding the six bits in flag1
assign {flag2}=flag1+A[6]+B[6];	//calculating the sum of flag1 and the 7th bit of A and B and storing the carry generated by the sum in flag2 (flag2 is used for parity)

//This block subtracts  A and B and stores the carry in carry2 
assign c1=~B+8'b00000001;		//flipping the bits and adding one(to make B as 2's complemented number)
assign {carry2,a2}=A[7:0]+c1[7:0];		//this logic is same as that of addition
assign {flag3}=A[5:0]+c1[5:0];
assign {flag4}=flag3+A[6]+c1[6];

assign a4=A&B;
assign a5=A|B;
assign a6=A^B;
assign a7=~B;
assign a22=A<<B;
assign a23=A>>B;

//this code will do arithmeric right shift
assign a24 = B[3:0] == 4'b0000 ?A:(B[3:0] == 4'b0001 ?{A[7],A[7],A[6:1]}:(B[3:0] == 4'b0010 ?{A[7],A[7],A[7],A[6:2]}:(B[3:0] == 4'b0011 ?{A[7],A[7],A[7],A[7],A[6:3]}:(B[3:0] == 4'b0100 ?{A[7],A[7],A[7],A[7],A[7],A[6:4]}:(B[3:0] == 4'b0101 ?{A[7],A[7],A[7],A[7],A[7],A[7],A[6:5]}:(B[3:0] == 4'b0110 ?{A[7],A[7],A[7],A[7],A[7],A[7],A[7],A[6]}:{A[7],A[7],A[7],A[7],A[7],A[7],A[7],A[7]})))))); 

//this code will assign the value to ans_temp according to opcode(ans_temp is the value which ans_ex will get)
assign ans_temp = (op_dec==5'b00000 ?a1:(op_dec==5'b00001 ?a2:(op_dec==5'b00010 ?B:(op_dec==5'b00100 ?a4:(op_dec==5'b00101 ?a5:(op_dec==5'b00110 ?a6:(op_dec==5'b00111 ?a7:(op_dec==5'b01000 ?a1:(op_dec==5'b01001 ?a2:(op_dec==5'b01010 ?B:(op_dec==5'b01100 ?a4:(op_dec==5'b01101 ?a5:(op_dec==5'b01110 ?a6:(op_dec==5'b01111 ?a7:(op_dec==5'b10000 ?ans_ex:(op_dec==5'b10001 ?ans_ex:(op_dec==5'b10100 ?A:(op_dec==5'b10101 ?A:(op_dec==5'b10110 ?data_in:(op_dec==5'b10111 ?ans_ex:(op_dec==5'b11000 ?ans_ex:(op_dec==5'b11001 ?a22:(op_dec==5'b11010 ?a23:(op_dec==5'b11011 ?a24:(op_dec==5'b11100 ?ans_ex:(op_dec==5'b11101 ?ans_ex:(op_dec==5'b11110 ?ans_ex:(op_dec==5'b11111 ?ans_ex:8'b00000000))))))))))))))))))))))))))));

//storing the bits of flag in r1,r2,r3,r4 using flip flops
d_flipflop dff1(flag_ex[0],r1,reset,clk);
d_flipflop dff2(flag_ex[1],r2,reset,clk);
d_flipflop dff3(flag_ex[2],r3,reset,clk);
d_flipflop dff4(flag_ex[3],r4,reset,clk);

//This assign 
assign flag_temp = (op_dec==5'b00000) ?flag2:(op_dec==5'b00001 ?flag4:(op_dec==5'b01000 ?flag2:(op_dec==5'b01001 ?flag4:1'b0)));

//the assignment statement from t1 to t6 are for grouping the opcodes which affect similar flag

assign t1 = (op_dec==5'b00000 || op_dec==5'b00001 || op_dec==5'b01000 || op_dec==5'b01001);

assign t2 = (op_dec==5'b00010 || op_dec==5'b00100 || op_dec==5'b00101 || op_dec==5'b00110 || op_dec==5'b00111 || op_dec==5'b01010 || op_dec==5'b01100 || op_dec==5'b01101 || op_dec==5'b01110 || op_dec==5'b01111 || op_dec==5'b10110 || op_dec==5'b11001 || op_dec==5'b11010 || op_dec==5'b11011);

assign t3 = (op_dec==5'b10000 || op_dec==5'b10001);

assign t4 = (op_dec==5'b10100 || op_dec==5'b10101 || op_dec==5'b10111 || op_dec==5'b11000 || op_dec==5'b11100 || op_dec==5'b11101 || op_dec==5'b11110 || op_dec==5'b11111);

assign carry = (op_dec == 5'b00000 ? carry1:(op_dec == 5'b00001 ? carry2:(op_dec == 5'b01000 ? carry1:(op_dec == 5'b01001 ? carry2:1'b0))));

//t5 calculates the value of zero flag by oring all the bits of ans_temp 
assign t5 = ~(ans_temp[7] | ans_temp[6] | ans_temp[5] | ans_temp[4] | ans_temp[3] | ans_temp[2] | ans_temp[1] | ans_temp[0]);

//t6 calculates the value of parity flag by xoring all the bits of ans_temp 
assign t6 = (ans_temp[7]^ans_temp[6]^ans_temp[5]^ans_temp[4]^ans_temp[3]^ans_temp[2]^ans_temp[1]^ans_temp[0]);


//assigning the value of flag_ex according to the opcodes
assign flag_ex[0] = (t1==1 ? carry :(t2==1 ?1'b0:(t3==1 ?1'b0:(t4==1 ?r1:1'b0))));

assign flag_ex[1] = (t1==1 ? t5 :(t2==1 ?t5:(t3==1 ?1'b0:(t4==1 ?r2:1'b0))));

assign flag_ex[2] = (t1==1 ?flag_ex[0]^flag_temp:(t2==1 ?1'b0:(t3==1 ?1'b0:(t4==1 ?r3:1'b0))));

assign flag_ex[3] = (t1==1 ? t6 :(t2==1 ?t6:(t3==1 ?1'b0:(t4==1 ?r4:1'b0))));

//assigning the value to data_out_buff
assign data_out_buff = (op_dec == 5'b10111) ? A:data_out;

assign ans_ex_t = (reset==1'b1) ?ans_temp :8'b00000000;		//ans_ex_t is a temporary wire that stores the value of ans_temp if reset is 1 otherwise it stores 8'b00000000 (ans_ex_t is a wire that gives the value to ans_ex at posedge clock)
assign data_out_t = (reset==1'b1) ? data_out_buff :8'b00000000;	//data_out_t is a temporary wire that stores the value of data_out_buff if reset is 1 otherwise it stores 8'b00000000 (data_out_t is a wire that gives the value to data_out at posedge clock)
assign B_Bypass_t = (reset==1'b1) ? B :8'b00000000;		//B_Bypass_t is a temporary wire that stores the value of B if reset is 1 otherwise it stores 8'b00000000 (B_Bypass_t is a wire that gives the value to B_Bypass at posedge clock)
assign mem_en_ex_t = (reset==1'b1) ?mem_en_dec :1'b0;		//mem_en_ex_t  is a temporary wire that stores the value of mem_en_dec if reset is 1 otherwise it stores 1'b0 (mem_en_ex_t  is a wire that gives the value to mem_en_ex at posedge clock)
assign mem_rw_ex_t = (reset==1'b1) ?mem_rw_dec :1'b0;		//mem_rw_ex_t  is a temporary wire that stores the value of mem_rw_dec if reset is 1 otherwise it stores 1'b0 (mem_rw_ex_t  is a wire that gives the value to mem_rw_ex at posedge clock)
assign mem_mux_sel_ex_t = (reset==1'b1) ?mem_mux_sel_dec :1'b0;	//mem_mux_sel_ex_t is a temporary wire that stores the value of mem_mux_sel_dec if reset is 1 otherwise it stores 1'b0 (mem_mux_sel_ex_t is a wire that gives the value to mem_mux_sel_ex at posedge clock)
assign RW_ex_t = (reset==1'b1) ?RW_dec :5'b00000;	//RW_ex_t is a temporary wire that stores the value of RW_dec if reset is 1 otherwise it stores 5'b00000 (RW_ex_t is a wire that gives the value to RW_ex at posedge clock)

always@(posedge clk) 
begin 
	RW_ex <= RW_ex_t;		//assigning the value of RW_ex_t to RW_ex at posedge clk
	mem_rw_ex <= mem_rw_ex_t;	//assigning the value of mem_rw_ex_t to mem_rw_ex at posedge clk
	mem_mux_sel_ex <= mem_mux_sel_ex_t; 	//assigning the value of mem_mux_sel_ex_t to mem_mux_sel_ex at posedge clk
	mem_en_ex <= mem_en_ex_t;		//assigning the value of mem_en_ex_t to mem_en_ex at posedge clk
	B_Bypass <= B_Bypass_t;		//assigning the value of B_Bypass_t to B_Bypass at posedge clk
	data_out <= data_out_t;		//assigning the value of data_out_t to data_out at posedge clk
	ans_ex <= ans_ex_t;	//assigning the value of ans_ex_t to ans_ex at posedge clk
end

endmodule
